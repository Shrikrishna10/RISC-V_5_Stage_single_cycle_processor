module mux_2_tb(input [31:0] d0, d1, input s, output y);

endmodule
