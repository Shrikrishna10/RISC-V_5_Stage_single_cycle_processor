module ifstage(input logic [31:0] 
