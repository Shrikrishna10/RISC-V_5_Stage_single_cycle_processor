module regis32(input logic [31:0] j,k, input clk, output logic [31:0] q, qn);

