module decoder(input [31:0]din, output [31:0] dout);

